module fast_test(
    input  [15:0] x0,
    input  [15:0] x1,
    input  [15:0] x2,
    input  [15:0] x3,
    input  [15:0] x4,
    input  [15:0] x5,
    input  [15:0] x6,
    input  [15:0] x7,
    output  [15:0] y0,
    output  [15:0] y1,
    output  [15:0] y2,
    output  [15:0] y3,
    output  [15:0] y4,
    output  [15:0] y5,
    output  [15:0] y6,
    output  [15:0] y7
);
// C1 = 0.49
// C2 = 0.46
// C3 = 0.42
// C4 = 0.35
// C5 = 0.28
// C6 = 0.19
// C7 = 0.10

// reg [20:0] X0 = {7'b0000000,x0,6'b000000};
// reg [20:0] X1 = {7'b0000000,x1,6'b000000};
// reg [20:0] X2 = {7'b0000000,x2,6'b000000};
// reg [20:0] X3 = {7'b0000000,x3,6'b000000};
// reg [20:0] X4 = {7'b0000000,x4,6'b000000};
// reg [20:0] X5 = {7'b0000000,x5,6'b000000};
// reg [20:0] X6 = {7'b0000000,x6,6'b000000};
// reg [20:0] X7 = {7'b0000000,x7,6'b000000};

reg [25:0] C1 = 25'b0000000000000000_0111110101;
reg [25:0] C2 = 25'b0000000000000000_0111010111;
reg [25:0] C3 = 25'b0000000000000000_0110101110;
reg [25:0] C4 = 25'b0000000000000000_0101100110; 
reg [25:0] C5 = 25'b0000000000000000_0100011110;
reg [25:0] C6 = 25'b0000000000000000_0011000010;
reg [25:0] C7 = 25'b0000000000000000_0001100110;
//------------------------------------------------------------------------------------------------
reg [25:0] s07;
reg [25:0] s16;
reg [25:0] s25;
reg [25:0] s34;
reg [25:0] temp1;
reg [25:0] temp2;
reg [25:0] s07341625;
reg [25:0] Y0;

qadd #(10,26) u1(.a({x0,10'b0000000000}),.b({x7,10'b0000000000}),.c(s07));
qadd #(10,26) u2(.a({x1,10'b0000000000}),.b({x6,10'b0000000000}),.c(s16));
qadd #(10,26) u3(.a({x2,10'b0000000000}),.b({x5,10'b0000000000}),.c(s25));
qadd #(10,26) u4(.a({x3,10'b0000000000}),.b({x4,10'b0000000000}),.c(s34));
qadd #(10,26) u5(.a(s07),.b(s16),.c(temp1));
qadd #(10,26) u6(.a(s25),.b(s34),.c(temp2));
qadd #(10,26) u7(.a(temp1),.b(temp2),.c(s07341625));
qmult #(10,26) r1(.i_multiplicand(s07341625),.i_multiplier(C4),.o_result(Y0));
//-------------------------------------------------------------------------------------------------
reg [25:0] f0_7;
reg [25:0] f1_6;
reg [25:0] f2_5;
reg [25:0] f3_4;
reg [25:0] temp3;
reg [25:0] temp4;
reg [25:0] temp5;
reg [25:0] temp6;
reg [25:0] temp7;
reg [25:0] temp8;
reg [25:0] Y1;

qadd #(10,26) u8(.a({x0,10'b0000000000}),.b({~x7[15],x7[14:0],10'b0000000000}),.c(f0_7));
qadd #(10,26) u9(.a({x1,10'b0000000000}),.b({~x6[15],x6[14:0],10'b0000000000}),.c(f1_6));
qadd #(10,26) u10(.a({x2,10'b0000000000}),.b({~x5[15],x5[14:0],10'b0000000000}),.c(f2_5));
qadd #(10,26) u11(.a({x3,10'b0000000000}),.b({~x4[15],x4[14:0],10'b0000000000}),.c(f3_4));
qmult #(10,26) r2(.i_multiplicand(f0_7),.i_multiplier(C1),.o_result(temp3));
qmult #(10,26) r3(.i_multiplicand(f1_6),.i_multiplier(C3),.o_result(temp4));
qmult #(10,26) r4(.i_multiplicand(f2_5),.i_multiplier(C5),.o_result(temp5));
qmult #(10,26) r5(.i_multiplicand(f3_4),.i_multiplier(C7),.o_result(temp6));
qadd #(10,26) u12(.a(temp3),.b(temp4),.c(temp7));
qadd #(10,26) u13(.a(temp5),.b(temp6),.c(temp8));
qadd #(10,26) u14(.a(temp7),.b(temp8),.c(Y1));
//-------------------------------------------------------------------------------------------------
reg [25:0] s07_34;
reg [25:0] s16_25;
reg [25:0] temp9;
reg [25:0] temp10;
reg [25:0] Y2;
qadd #(10,26) u15(.a(s07),.b({(~s34[25]),s34[24:0]}),.c(s07_34));
qadd #(10,26) u16(.a(s16),.b({(~s25[25]),s25[24:0]}),.c(s16_25));
qmult #(10,26) r6(.i_multiplicand(s07_34),.i_multiplier(C2),.o_result(temp9));
qmult #(10,26) r7(.i_multiplicand(s16_25),.i_multiplier(C6),.o_result(temp10));
qadd #(10,26) u17(.a(temp9),.b(temp10),.c(Y2));
//--------------------------------------------------------------------------------------------------
reg [25:0] f0_7_C3;
reg [25:0] f1_6_C7;
reg [25:0] f2_5_C1;
reg [25:0] f3_4_C5;
reg [25:0] temp11;
reg [25:0] temp12;
reg [25:0] Y3;

qmult #(10,26) r8(.i_multiplicand(f0_7),.i_multiplier(C3),.o_result(f0_7_C3));
qmult #(10,26) r9(.i_multiplicand(f1_6),.i_multiplier({~C7[25],C7[24:0]}),.o_result(f1_6_C7));
qmult #(10,26) r10(.i_multiplicand(f2_5),.i_multiplier({~C1[25],C1[24:0]}),.o_result(f2_5_C1));
qmult #(10,26) r11(.i_multiplicand(f3_4),.i_multiplier({~C5[25],C5[24:0]}),.o_result(f3_4_C5));
qadd #(10,26) u18(.a(f0_7_C3),.b(f1_6_C7),.c(temp11));
qadd #(10,26) u19(.a(f2_5_C1),.b(f3_4_C5),.c(temp12));
qadd #(10,26) u20(.a(temp11),.b(temp12),.c(Y3));
//-----------------------------------------------------------------------------------------------------
reg [25:0] s0734;
reg [25:0] s0734_16;
reg [25:0] s0734_16_25;
reg [25:0] Y4;
qadd #(10,26) u21(.a(s07),.b(s34),.c(s0734));
qadd #(10,26) u22(.a(s0734),.b({~s16[25],s16[24:0]}),.c(s0734_16));
qadd #(10,26) u23(.a(s0734_16),.b({~s25[25],s25[24:0]}),.c(s0734_16_25));
qmult #(10,26) r12(.i_multiplicand(s0734_16_25),.i_multiplier(C4),.o_result(Y4));
//------------------------------------------------------------------------------------------------------
reg [25:0] f0_7_C5;
reg [25:0] f1_6_C1;
reg [25:0] f2_5_C7;
reg [25:0] f3_4_C3;
reg [25:0] temp13;
reg [25:0] temp14;
reg [25:0] Y5;
qmult #(10,26) r13(.i_multiplicand(f0_7),.i_multiplier(C5),.o_result(f0_7_C5));
qmult #(10,26) r14(.i_multiplicand(f1_6),.i_multiplier({~C1[25],C1[24:0]}),.o_result(f1_6_C1));
qmult #(10,26) r15(.i_multiplicand(f2_5),.i_multiplier(C7),.o_result(f2_5_C7));
qmult #(10,26) r16(.i_multiplicand(f3_4),.i_multiplier(C3),.o_result(f3_4_C3));
qadd #(10,26) u24(.a(f0_7_C5),.b(f1_6_C1),.c(temp13));
qadd #(10,26) u25(.a(f2_5_C7),.b(f3_4_C3),.c(temp14));
qadd #(10,26) u26(.a(temp13),.b(temp14),.c(Y5));
//-------------------------------------------------------------------------------------------------------
reg [25:0] s07_34_C6;
reg [25:0] s16_25_C2;
reg [25:0] Y6;
qmult #(10,26) r17(.i_multiplicand(s07_34),.i_multiplier(C6),.o_result(s07_34_C6));
qmult #(10,26) r18(.i_multiplicand(s16_25),.i_multiplier({~C2[25],C2[24:0]}),.o_result(s16_25_C2));
qadd #(10,26) u27(.a(s07_34_C6),.b(s16_25_C2),.c(Y6));
//--------------------------------------------------------------------------------------------------------
reg [25:0] f0_7_C7;
reg [25:0] f1_6_C5;
reg [25:0] f2_5_C3;
reg [25:0] f3_4_C1;
reg [25:0] temp15;
reg [25:0] temp16;
reg [25:0] Y7;
qmult #(10,26) r19(.i_multiplicand(f0_7),.i_multiplier(C7),.o_result(f0_7_C7));
qmult #(10,26) r20(.i_multiplicand(f1_6),.i_multiplier({~C5[25],C5[24:0]}),.o_result(f1_6_C5));
qmult #(10,26) r21(.i_multiplicand(f2_5),.i_multiplier(C3),.o_result(f2_5_C3));
qmult #(10,26) r22(.i_multiplicand(f3_4),.i_multiplier({~C1[25],C1[24:0]}),.o_result(f3_4_C1));
qadd #(10,26) u28(.a(f0_7_C7),.b(f1_6_C5),.c(temp15));
qadd #(10,26) u29(.a(f2_5_C3),.b(f3_4_C1),.c(temp16));
qadd #(10,26) u30(.a(temp15),.b(temp16),.c(Y7));
//---------------------------------------------------------------------------------------------------------



always_comb begin
    y0 = Y0[25:10];
    y1 = Y1[25:10];
    y2 = Y2[25:10];
    y3 = Y3[25:10];
    y4 = Y4[25:10];
    y5 = Y5[25:10];
    y6 = Y6[25:10];
    y7 = Y7[25:10];

end




endmodule




