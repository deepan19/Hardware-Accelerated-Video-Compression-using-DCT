module fast_test(
    input  [14:0] x0,
    input  [14:0] x1,
    input  [14:0] x2,
    input  [14:0] x3,
    input  [14:0] x4,
    input  [14:0] x5,
    input  [14:0] x6,
    input  [14:0] x7,
    output  [14:0] y0,
    output  [14:0] y1,
    output  [14:0] y2,
    output  [14:0] y3,
    output  [14:0] y4,
    output  [14:0] y5,
    output  [14:0] y6,
    output  [14:0] y7
);
// C1 = 0.49
// C2 = 0.46
// C3 = 0.42
// C4 = 0.35
// C5 = 0.28
// C6 = 0.19
// C7 = 0.10

// reg [20:0] X0 = {7'b0000000,x0,6'b000000};
// reg [20:0] X1 = {7'b0000000,x1,6'b000000};
// reg [20:0] X2 = {7'b0000000,x2,6'b000000};
// reg [20:0] X3 = {7'b0000000,x3,6'b000000};
// reg [20:0] X4 = {7'b0000000,x4,6'b000000};
// reg [20:0] X5 = {7'b0000000,x5,6'b000000};
// reg [20:0] X6 = {7'b0000000,x6,6'b000000};
// reg [20:0] X7 = {7'b0000000,x7,6'b000000};

reg [24:0] C1 = 24'b000000000000000_0111110101;
reg [24:0] C2 = 24'b000000000000000_0111010111;
reg [24:0] C3 = 24'b000000000000000_0110101110;
reg [24:0] C4 = 24'b000000000000000_0101100110; 
reg [24:0] C5 = 24'b000000000000000_0100011110;
reg [24:0] C6 = 24'b000000000000000_0011000010;
reg [24:0] C7 = 24'b000000000000000_0001100110;
//------------------------------------------------------------------------------------------------
reg [24:0] s07;
reg [24:0] s16;
reg [24:0] s25;
reg [24:0] s34;
reg [24:0] temp1;
reg [24:0] temp2;
reg [24:0] s07341625;
reg [24:0] Y0;

qadd #(10,25) u1(.a({x0,10'b0000000000}),.b({x7,10'b0000000000}),.c(s07));
qadd #(10,25) u2(.a({x1,10'b0000000000}),.b({x6,10'b0000000000}),.c(s16));
qadd #(10,25) u3(.a({x2,10'b0000000000}),.b({x5,10'b0000000000}),.c(s25));
qadd #(10,25) u4(.a({x3,10'b0000000000}),.b({x4,10'b0000000000}),.c(s34));
qadd #(10,25) u5(.a(s07),.b(s16),.c(temp1));
qadd #(10,25) u6(.a(s25),.b(s34),.c(temp2));
qadd #(10,25) u7(.a(temp1),.b(temp2),.c(s07341625));
qmult #(10,25) r1(.i_multiplicand(s07341625),.i_multiplier(C4),.o_result(Y0));
//-------------------------------------------------------------------------------------------------
reg [24:0] f0_7;
reg [24:0] f1_6;
reg [24:0] f2_5;
reg [24:0] f3_4;
reg [24:0] temp3;
reg [24:0] temp4;
reg [24:0] temp5;
reg [24:0] temp6;
reg [24:0] temp7;
reg [24:0] temp8;
reg [24:0] Y1;

qadd #(10,25) u8(.a({x0,10'b0000000000}),.b({~x7[14],x7[13:0],10'b0000000000}),.c(f0_7));
qadd #(10,25) u9(.a({x1,10'b0000000000}),.b({~x6[14],x6[13:0],10'b0000000000}),.c(f1_6));
qadd #(10,25) u10(.a({x2,10'b0000000000}),.b({~x5[14],x5[13:0],10'b0000000000}),.c(f2_5));
qadd #(10,25) u11(.a({x3,10'b0000000000}),.b({~x4[14],x4[13:0],10'b0000000000}),.c(f3_4));
qmult #(10,25) r2(.i_multiplicand(f0_7),.i_multiplier(C1),.o_result(temp3));
qmult #(10,25) r3(.i_multiplicand(f1_6),.i_multiplier(C3),.o_result(temp4));
qmult #(10,25) r4(.i_multiplicand(f2_5),.i_multiplier(C5),.o_result(temp5));
qmult #(10,25) r5(.i_multiplicand(f3_4),.i_multiplier(C7),.o_result(temp6));
qadd #(10,25) u12(.a(temp3),.b(temp4),.c(temp7));
qadd #(10,25) u13(.a(temp5),.b(temp6),.c(temp8));
qadd #(10,25) u14(.a(temp7),.b(temp8),.c(Y1));
//-------------------------------------------------------------------------------------------------
reg [24:0] s07_34;
reg [24:0] s16_25;
reg [24:0] temp9;
reg [24:0] temp10;
reg [24:0] Y2;
qadd #(10,25) u15(.a(s07),.b({(~s34[24]),s34[23:0]}),.c(s07_34));
qadd #(10,25) u16(.a(s16),.b({(~s25[24]),s25[23:0]}),.c(s16_25));
qmult #(10,25) r6(.i_multiplicand(s07_34),.i_multiplier(C2),.o_result(temp9));
qmult #(10,25) r7(.i_multiplicand(s16_25),.i_multiplier(C6),.o_result(temp10));
qadd #(10,25) u17(.a(temp9),.b(temp10),.c(Y2));
//--------------------------------------------------------------------------------------------------
reg [24:0] f0_7_C3;
reg [24:0] f1_6_C7;
reg [24:0] f2_5_C1;
reg [24:0] f3_4_C5;
reg [24:0] temp11;
reg [24:0] temp12;
reg [24:0] Y3;

qmult #(10,25) r8(.i_multiplicand(f0_7),.i_multiplier(C3),.o_result(f0_7_C3));
qmult #(10,25) r9(.i_multiplicand(f1_6),.i_multiplier({~C7[24],C7[23:0]}),.o_result(f1_6_C7));
qmult #(10,25) r10(.i_multiplicand(f2_5),.i_multiplier({~C1[24],C1[23:0]}),.o_result(f2_5_C1));
qmult #(10,25) r11(.i_multiplicand(f3_4),.i_multiplier({~C5[24],C5[23:0]}),.o_result(f3_4_C5));
qadd #(10,25) u18(.a(f0_7_C3),.b(f1_6_C7),.c(temp11));
qadd #(10,25) u19(.a(f2_5_C1),.b(f3_4_C5),.c(temp12));
qadd #(10,25) u20(.a(temp11),.b(temp12),.c(Y3));
//-----------------------------------------------------------------------------------------------------
reg [24:0] s0734;
reg [24:0] s0734_16;
reg [24:0] s0734_16_25;
reg [24:0] Y4;
qadd #(10,25) u21(.a(s07),.b(s34),.c(s0734));
qadd #(10,25) u22(.a(s0734),.b({~s16[24],s16[23:0]}),.c(s0734_16));
qadd #(10,25) u23(.a(s0734_16),.b({~s25[24],s25[23:0]}),.c(s0734_16_25));
qmult #(10,25) r12(.i_multiplicand(s0734_16_25),.i_multiplier(C4),.o_result(Y4));
//------------------------------------------------------------------------------------------------------
reg [24:0] f0_7_C5;
reg [24:0] f1_6_C1;
reg [24:0] f2_5_C7;
reg [24:0] f3_4_C3;
reg [24:0] temp13;
reg [24:0] temp14;
reg [24:0] Y5;
qmult #(10,25) r13(.i_multiplicand(f0_7),.i_multiplier(C5),.o_result(f0_7_C5));
qmult #(10,25) r14(.i_multiplicand(f1_6),.i_multiplier({~C1[24],C1[23:0]}),.o_result(f1_6_C1));
qmult #(10,25) r15(.i_multiplicand(f2_5),.i_multiplier(C7),.o_result(f2_5_C7));
qmult #(10,25) r16(.i_multiplicand(f3_4),.i_multiplier(C3),.o_result(f3_4_C3));
qadd #(10,25) u24(.a(f0_7_C5),.b(f1_6_C1),.c(temp13));
qadd #(10,25) u25(.a(f2_5_C7),.b(f3_4_C3),.c(temp14));
qadd #(10,25) u26(.a(temp13),.b(temp14),.c(Y5));
//-------------------------------------------------------------------------------------------------------
reg [24:0] s07_34_C6;
reg [24:0] s16_25_C2;
reg [24:0] Y6;
qmult #(10,25) r17(.i_multiplicand(s07_34),.i_multiplier(C6),.o_result(s07_34_C6));
qmult #(10,25) r18(.i_multiplicand(s16_25),.i_multiplier({~C2[24],C2[23:0]}),.o_result(s16_25_C2));
qadd #(10,25) u27(.a(s07_34_C6),.b(s16_25_C2),.c(Y6));
//--------------------------------------------------------------------------------------------------------
reg [24:0] f0_7_C7;
reg [24:0] f1_6_C5;
reg [24:0] f2_5_C3;
reg [24:0] f3_4_C1;
reg [24:0] temp15;
reg [24:0] temp16;
reg [24:0] Y7;
qmult #(10,25) r19(.i_multiplicand(f0_7),.i_multiplier(C7),.o_result(f0_7_C7));
qmult #(10,25) r20(.i_multiplicand(f1_6),.i_multiplier({~C5[24],C5[23:0]}),.o_result(f1_6_C5));
qmult #(10,25) r21(.i_multiplicand(f2_5),.i_multiplier(C3),.o_result(f2_5_C3));
qmult #(10,25) r22(.i_multiplicand(f3_4),.i_multiplier({~C1[24],C1[23:0]}),.o_result(f3_4_C1));
qadd #(10,25) u28(.a(f0_7_C7),.b(f1_6_C5),.c(temp15));
qadd #(10,25) u29(.a(f2_5_C3),.b(f3_4_C1),.c(temp16));
qadd #(10,25) u30(.a(temp15),.b(temp16),.c(Y7));
//---------------------------------------------------------------------------------------------------------



always_comb begin
    y0 = Y0[24:10];
    y1 = Y1[24:10];
    y2 = Y2[24:10];
    y3 = Y3[24:10];
    y4 = Y4[24:10];
    y5 = Y5[24:10];
    y6 = Y6[24:10];
    y7 = Y7[24:10];

end




endmodule




